(* Coq module loading the different ML components of the plugin *)

Declare ML Module "coqine_plugin".
